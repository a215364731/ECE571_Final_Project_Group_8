// Read ONLY, no rd enable needed. Read will be combinational
module imem(
    input logic [31:0] addr,
    output logic [31:0] data
);

endmodule