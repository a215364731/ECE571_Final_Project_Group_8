module riscv_core(
    input clk, reset_n
);

endmodule