module top_tb;

    logic clk, reset_n;

    riscv_core riscv_core(.*);

    initial begin
        
    end

endmodule